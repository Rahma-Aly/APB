import uvm_pkg::*;
`include "uvm_macros.svh"
import apb_pkg::*;

module hvl_top();

initial begin
	run_test("test");
end

endmodule: hvl_top
